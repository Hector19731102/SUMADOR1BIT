module C_XOR (A,B,OUT);
  input A;
  input B;
  output OUT;
  assign OUT=A^B;
endmodule
